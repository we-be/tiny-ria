module main

fn main() {
	println('Hello Charles Schwab!')
}
